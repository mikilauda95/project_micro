package CONSTANTS is
	constant IVDELAY : time := 0.1 ns;
	constant NDDELAY : time := 0.2 ns;
	constant NRDELAY : time := 0.2 ns;
	constant numbit : integer := 32;
	constant tp_mux: time := 3 ns;
	constant n : integer := 3;
	constant DRFAS: time := 0 ns ;
	constant DRFAC : time := 0 ns ;
end CONSTANTS;
