library ieee;
use ieee.std_logic_1164.all;
use work.log.all;

package types is

--	constant n_bit : natural := 16;
--	constant n_block : natural := 4;
--	constant log_n_bit : natural := log2_unsigned(n_bit);
--	constant log_n_block : natural := log2_unsigned(n_block);
--  type tree_conn is array (log_n_bit downto 0) of std_logic_vector((2*n_bit) downto 1);

end types;
